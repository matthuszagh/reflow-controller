.title KiCad schematic
R1 /D+ Net-_J1-Pad3_ 22
R2 Net-_J1-Pad2_ /D- 22
C6 VCC GND 1u
Y1 Net-_C4-Pad1_ Net-_C5-Pad1_ 8MHz
C4 Net-_C4-Pad1_ GND 26p
C5 Net-_C5-Pad1_ GND 26p
U1 GND Net-_C9-Pad2_ Net-_C9-Pad1_ VCC /SCK /SS /MISO MAX31855KASA
C3 GND VCC 0.1u
J2 Net-_C9-Pad2_ Net-_C9-Pad1_ Conn_01x02
J3 /MISO VCC /SCK /MOSI /RST GND Conn_02x03_Odd_Even
R3 VCC /RST 10k
D1 VCC /RST D
U2 /VBUS GND /VBUS NC_01 VCC AP2127K-3.3
C1 /VBUS GND 10u
C2 VCC GND 1u
Q1 Net-_Q1-Pad1_ GND Net-_J4-Pad2_ BC817
J4 VCC Net-_J4-Pad2_ Conn_01x02
J5 /RX /TX /VBUS GND Conn_01x04
C7 VCC GND 0.1u
C8 VCC GND 0.1u
U3 Net-_C4-Pad1_ Net-_C5-Pad1_ GND VCC NC_02 NC_03 NC_04 /RX /TX NC_05 NC_06 NC_07 NC_08 /SS /SCK /MOSI /MISO NC_09 NC_10 NC_11 NC_12 NC_13 /RELAY /RST NC_14 NC_15 VCC GND /D+ /D- VCC VCC ATmega8U2-AU
J1 /VBUS Net-_J1-Pad2_ Net-_J1-Pad3_ NC_16 GND GND USB_B_Mini
R6 Net-_Q1-Pad1_ /RELAY 1k
C9 Net-_C9-Pad1_ Net-_C9-Pad2_ 10n
R5 VCC /SS 10k
D2 GND Net-_D2-Pad2_ LED
R4 VCC Net-_D2-Pad2_ 240
.end
